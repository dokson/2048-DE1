LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
 
PACKAGE GAME_UTILS IS
	FUNCTION INT_TO7SEG (A:INTEGER) 
		RETURN STD_LOGIC_VECTOR;
END GAME_UTILS;
 
 
PACKAGE BODY GAME_UTILS IS
	
FUNCTION DIGIT_TO7SEG (A:INTEGER) RETURN STD_LOGIC_VECTOR IS
	
-- Risultato: uscita 7 bit per 7 segmenti
VARIABLE RESULT: STD_LOGIC_VECTOR(6 downto 0);

BEGIN
	CASE A IS
		WHEN 0 => RESULT:="1000000";
		WHEN 1 => RESULT:="1111001";
		WHEN 2 => RESULT:="0100100";
		WHEN 3 => RESULT:="0110000";
		WHEN 4 => RESULT:="0011001";
		WHEN 5 => RESULT:="0010010";
		WHEN 6 => RESULT:="0000010";
		WHEN 7 => RESULT:="1111000";
		WHEN 8 => RESULT:="0000000";
		WHEN 9 => RESULT:="0010000";
		WHEN OTHERS => RESULT:=(OTHERS=>'0');
	END CASE;
	RETURN RESULT;

END DIGIT_TO7SEG;
END GAME_UTILS;