LIBRARY IEEE;
use IEEE.STD_LOGIC_1164.ALL;

PACKAGE GAME_TYPES IS
	
	type GAME_GRID is array (3 downto 0, 3 downto 0) of integer;

END GAME_TYPES;
