LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE WORK.GAME_TYPES.ALL;
USE WORK.GAME_UTILS.ALL;

entity GAME_BOX is
	generic
	(
		XPOS 	: in NATURAL;
		YPOS 	: in NATURAL
	);
	port
	(
		-- INPUT
		clk		: IN STD_LOGIC;
		pixel_x : IN INTEGER RANGE 0 to 1000;
		pixel_y : IN INTEGER RANGE 0 to 500;
		number	: IN INTEGER RANGE 0 to 2500; 		
		
		-- OUTPUT
		color	: OUT STD_LOGIC_VECTOR(11 downto 0); -- colore attuale del box
		drawBox : OUT STD_LOGIC := '0' 	-- disegna il box quando drawBox = 1
	);
end GAME_BOX;

architecture box_arch of GAME_BOX is
	-- Dimensioni fisse di tutti i box
	constant larghezza 	: integer := 150; 	
	constant altezza 	: integer := 105;
	-- Coordinate finali del cubo sullo schermo
	constant MAX_X 		: integer := XPOS + larghezza; -- larghezza
	constant MAX_Y 		: integer := YPOS + altezza; -- altezza
	-- Coordinate delle cifre sullo schermo
	constant X_CHAR		: integer := XPOS + larghezza/2;
	constant Y_CHAR		: integer := YPOS + altezza/2;
	 
	-- Segnali per la scrittura dei numeri a video
	signal numberToDraw1: character;
	signal numberToDraw2: character;
	signal numberToDraw3: character;
	signal numberToDraw4: character;
	signal drawNum1		: std_logic;
	signal drawNum2		: std_logic;
	signal drawNum3		: std_logic;
	signal drawNum4		: std_logic;

begin
	CH1: entity work.GAME_CHDISPLAY
	generic map
	(
		XPOS => X_CHAR-20,
		YPOS => Y_CHAR
	)
	port map
	(
		pixel_x 	=> pixel_x,
		pixel_y		=> pixel_y,
		char_code 	=> numberToDraw1,
		drawChar 	=> drawNum1
	);
	CH2: entity work.GAME_CHDISPLAY
	generic map
	(
		XPOS => X_CHAR-10,
		YPOS => Y_CHAR
	)
	port map
	(
		pixel_x		=> pixel_x,
		pixel_y		=> pixel_y,
		char_code 	=> numberToDraw2,
		drawChar 	=> drawNum2
	);
	CH3: entity work.GAME_CHDISPLAY
	generic map
	(
		XPOS => X_CHAR,
		YPOS => Y_CHAR
	)
	port map
	(
		pixel_x 	=> pixel_x,
		pixel_y		=> pixel_y,
		char_code 	=> numberToDraw3,
		drawChar 	=> drawNum3
	);
	CH4: entity work.GAME_CHDISPLAY
	generic map
	(
		XPOS => X_CHAR+10,
		YPOS => Y_CHAR
	)
	port map
	(
		pixel_x 	=> pixel_x,
		pixel_y		=> pixel_y,
		char_code 	=> numberToDraw4,
		drawChar 	=> drawNum4
	);
	
	valueChange : process(number, drawNum1, drawNum2, drawNum3, drawNum4, clk)
		variable digit4, digit3, digit2, digit1	: integer range 0 to 9;
	begin
		if(clk'event and clk = '1')
		then
			if not(drawNum1 = '1' or drawNum2 = '1' or drawNum3 = '1' or drawNum4 = '1')
			then
				case number is
					when 0 => 
						color <= COLOR_0;
					when 2 => 
						color <= COLOR_2;
					when 4 => 
						color <= COLOR_4;
					when 8 => 
						color <= COLOR_8;
					when 16 => 
						color <= COLOR_16;
					when 32 => 
						color <= COLOR_32;
					when 64 => 
						color <= COLOR_64;
					when 128 =>
						color <= COLOR_128;
					when 256 =>
						color <= COLOR_256;
					when 512 =>
						color <= COLOR_512;
					when 1024 =>
						color <= COLOR_1024;
					when 2048 =>
						color <= COLOR_2048;
					when others => 
						color <= COLOR_BLACK;
				end case;
				
				splitNumber(number, digit4, digit3, digit2, digit1);
				
				if(digit4 = 0)
				then
					numberToDraw1 <= NUL;
					if(digit3 = 0)
					then
						numberToDraw2 <= NUL;
						if(digit2 = 0)
						then
							numberToDraw3 <= NUL;
							if(digit1 = 0)
							then
								numberToDraw4 <= NUL;
							else
								numbertoDraw4 <= digit_to_char(digit1);
							end if;
						else
							numberToDraw3 <= digit_to_char(digit2);
							numberToDraw4 <= digit_to_char(digit1);
						end if;
					else
						numberToDraw2 <= digit_to_char(digit3);
						numberToDraw3 <= digit_to_char(digit2);
						numberToDraw4 <= digit_to_char(digit1);
					end if;
				else
					numberToDraw1 <= digit_to_char(digit4);
					numberToDraw2 <= digit_to_char(digit3);
					numberToDraw3 <= digit_to_char(digit2);
					numberToDraw4 <= digit_to_char(digit1);
				end if;
				
			else
				color <= COLOR_BLACK;
			end if;
		end if;
	end process valueChange;
	
	drawBox <= '1' 
	when 
		(pixel_x >= XPOS and pixel_x <= MAX_X and pixel_y >= YPOS and pixel_y <= MAX_Y)
	else
		'0';	
	
end box_arch;
